module bstone
