module bstone

struct Player {

}

fn (p Player) handle_packet(packet vraklib.Packet) {
    
}