module raknet

struct RakLib {

}